module sc_decoder(SC,Ti);

output [15:0] Ti;
input [3:0] SC;

reg [15:0] Ti;

always @ (SC)

	case(SC)
	 
 	4'b0000 : Ti = 16'b0000_0000_0001;
	4'b0001 : Ti = 16'b0000_0000_0010;
	4'b0010 : Ti = 16'b0000_0000_0100;
	4'b0011 : Ti = 16'b0000_0000_1000;
	4'b0100 : Ti = 16'b0000_0001_0000;
	4'b0101 : Ti = 16'b0000_0010_0000;
	4'b0110 : Ti = 16'b0000_0100_0000;
	4'b0111 : Ti = 16'b0000_1000_0000;
	
	default : Ti = 16'b0000_0000_0000;

	endcase

endmodule
